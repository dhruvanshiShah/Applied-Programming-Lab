There could be junk here!
Since this portion does not belong to circuit definition.
.circuit
V1 GND 1 dc 10    # There can be comment here
R1 1 2 1e3
R2 2 3 1e3
R3 3 4 1e3
R4 4 5 1e3      # comment can be in any line
R5 2 GND 2e3
R6 3 GND 2e3
R7 4 GND 2e3
R8 5 GND 2e3
.end
There could be junk here!
Since this portion does not belong to circuit definition.
